`timescale 1ns / 1ps



module id_ex(

    input   logic       clk,reset,
    input   logic [1:0] ResultSrcD,
    input   logic       MemWriteD,
    input   logic       ALUSrcD,
    input   logic       RegWriteD, JumpD,BranchD,
    input   logic [2:0] ALUControlD,
    

                        
    

    );
endmodule
